
`define  time_period       8
`define  ffi_max           3
`define  receptive_field   8
`define  neurons_per_layer 16

