`ifndef INTERNAL_DEFINES_VH_
`define INTERNAL_DEFINES_VH_

`define  time_period            16
`define  log_time_period	4
`define  testing_period         8
`define  ffi_max                5
`define  num_spikes             8
`define  log_num_spikes		3
`define  neurons_per_layer     16
`define  log_neurons_per_layer  4
`define  THRESHOLD              14
`define  WBITS                  3    
`define  wmax                   7
 
`endif /* INTERNAL_DEFINES_VH_ */
