
`define  time_period       8
`define  ffi_max           3
`define  num_spikes   8
`define  neurons_per_layer 16
`define  THRESHOLD         2
`define  WBITS             2    // num bits in weights
`define  wmax               7
