`ifndef INTERNAL_DEFINES_VH_
`define INTERNAL_DEFINES_VH_

`define  time_period       8
`define  ffi_max           3
`define  num_spikes    8
`define  neurons_per_layer 16
`define  THRESHOLD         2
`define  WBITS             3    
`define  wmax               7

`endif /* INTERNAL_DEFINES_VH_ */
